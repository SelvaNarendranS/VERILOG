module top_module(
    input clk,
    input areset,    // Asynchronous reset to state B
    input in,
    output out); 

    parameter A=0, B=1; 
    reg state, next_state;

    always @(*) begin    // This is a combinational always block
        next_state = 1'bx;
        
        case(state)
            B :if(in == 0)
                    next_state = A;
                else
                    next_state = B;
            A : if(in == 0)
                next_state = B;            
            else
                next_state = A;
        endcase
    end

    always @(posedge clk or posedge areset) begin    // This is a sequential always block
        if(areset)
            state <= B;
        else
            state <= next_state;
    end

    // Output logic
    assign out = (state == B);

endmodule
