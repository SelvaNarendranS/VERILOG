// Gate level implementation

module nand_gate( input a, b, output c);

  // assign c = ~(a & b);
  nand(c , a, b);
  
endmodule
