// // Gate level implementation

module or_gate(input a,b, output c);

	//assign c = a + b;
	or (c, a, b);

endmodule


