module top_module (
    input clk,
    input slowena,
    input reset,
    output [3:0] q);
    
    always @(posedge clk) begin
        if(reset)
            q <= 1'b0;
        else if(slowena) begin
            if(q > 8)
            	q <= 1'b0;
        	else 
            	q <= q + 1'b1;
        end
    end

endmodule
