// Gate level implementation

module not_gate(input a , output b );

	//assign b = ~a;
	not(b, a);

endmodule
